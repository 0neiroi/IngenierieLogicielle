�� sr projet.Jeu2048.model.Grille��H�� I scoreI 	valeurMaxL grillet Ljava/util/HashSet;xp       sr java.util.HashSet�D�����4  xpw   ?@     sr projet.Jeu2048.model.Case�-�ie�� Z fusionI valeurI xI yL maGrillet Lprojet/Jeu2048/model/Grille;xp       ����q ~ sq ~        ����q ~ x